library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;
library work;


entity ControlUnit is
	port(

	);
	
end ControlUnit;

architecture behaivour of ControlUnit is
begin


end behaivour;