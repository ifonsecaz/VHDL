-- Aquí vamos a hacer el proyecto final.