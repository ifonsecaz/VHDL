library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;


entity InstructionMemory is
	port(
		
	);
	
end InstructionMemory;

architecture behaivour of InstructionMemory is

begin


end behaivour;