library ieee;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all;

entity Practica5 is
	port
	(
		CLK : in std_logic;
		reset: in std_logic;
		write_sig : in std_logic;
		D_address : in std_logic_vector(2 downto 0);
		A_address : in std_logic_vector(2 downto 0);
		B_address : in std_logic_vector(2 downto 0);
		D_data    : in std_logic_vector(15 downto 0);
		A_data    : out std_logic_vector(15 downto 0);
		B_data    : out std_logic_vector(15 downto 0);
		disp_address :  in std_logic_Vector(2 downto 0);
		disp_out     : out std_logic_vector(15 downto 0);
		r0_debug  : out std_logic_vector(15 downto 0);
		r1_debug  : out std_logic_vector(15 downto 0);
		r2_debug  : out std_logic_vector(15 downto 0);
		r3_debug  : out std_logic_vector(15 downto 0);
		r4_debug  : out std_logic_vector(15 downto 0);
		r5_debug  : out std_logic_vector(15 downto 0);
		r6_debug  : out std_logic_vector(15 downto 0);
		r7_debug  : out std_logic_vector(15 downto 0));
end Practica5;


architecture behavior of Practica5 is
type mem_type is array (2**3 - 1 downto 0) of std_logic_vector(15 downto 0) ;
signal mem : mem_type := (others => X"0000"); --X"0000";

signal cte : std_logic_vector(15 downto 0);
--signal A_res : std_logic_vector(15 downto 0) : X"0000" ;
begin
	cte <= X"0002";
	process (CLK)
	begin
		if (CLK'event AND CLK = '1') then
			if RESET = '1' then
				mem <= (others => X"0000");
			elsif write_sig = '1' then
				mem(to_integer(unsigned(D_address))) <= D_data;
			end if;
			
			
			
		end if;
	end process;
	A_data <= mem(to_integer(unsigned(A_address)));
			B_data <= mem(to_integer(unsigned(B_address)));
			disp_out <= mem(to_integer(unsigned(disp_address)));
			--mem(to_integer(unsigned(cte))) <= X"9876";
			r0_debug <= mem(0);
			r1_debug <= mem(1);
			r2_debug <= mem(2);
			r3_debug <= mem(3);
			r4_debug <= mem(4);
			r5_debug <= mem(5);
			r6_debug <= mem(6);
			r7_debug <= mem(7);
end behavior;
		