library ieee;

use ieee.std_logic_arith.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity CircuitoLogico is

	port(
				A : in std_logic_vector(0 to 15);
				B : in std_logic_vector(0 to 15);
				S : in std_logic_vector(0 to 1);
				G : out std_logic_vector(0 to 15));

end CircuitoLogico;


architecture behavior of CircuitoLogico is
	begin
		with S select
			G <=  A and B when "00",
					A or B when "01",
					A xor B when "10",
					not(A) when "11",
					"XXXXXXXXXXXXXXXX" when others;
end behavior;