library ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity CircuitoAritmetico is

	port(
			A    : IN STD_LOGIC_VECTOR(0 to 15);
			B    : IN STD_LOGIC_VECTOR(0 to 15);
			S    : IN STD_LOGIC_VECTOR(0 to 1);
			CIN  : IN STD_LOGIC;
			G    : OUT STD_LOGIC_VECTOR(0 to 15);
			COUT : OUT STD_LOGIC);
			
end CircuitoAritmetico;


architecture behavior of CircuitoAritmetico is
signal Y: STD_LOGIC_VECTOR(0 to 15) := "0000000000000000";
begin
	with S select
			Y <=  "0000000000000000" when "00",
					B                  when "01",
					not(B)             when "10",
					"1111111111111111" when "11",
					"XXXXXXXXXXXXXXXX" when others;
	G <= A + Y + CIN;
end behavior;